
interface spi_4wire_agent_if(input clk);
        
        logic ce ;
        logic sclk;
        logic sdi;
        logic sdo;


endinterface